`ifndef params
`define params

    parameter DEPTH         = 8;
    parameter CLK_PERIOD    = 10;
    
`endif